`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Jafet Chaves Barrantes
// 
// Create Date:    18:28:34 03/22/2016 
// Design Name: 
// Module Name:    Generador_Caracteres 
// Project Name: 
// Target Devices: 
// Tool versions: 
/* Description: Este m�dulo se encarga de generar el texto que se requiere en la imagen del monitor,
se compone de una memoria RAM (character_memory), una memoria ROM (font_rom)*/
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module generador_caracteres(
    );


endmodule
